------------------------------------------------------------------------------
--  File: func_one_tb.vhd
------------------------------------------------------------------------------
--Adder testbench
library IEEE;
use IEEE.std_logic_1164.all;

--Testbench entity is always empty
entity funcOneTestBench is
end funcOneTestBench;

architecture Bench of funcOneTestBench is 
	
begin
	

end Bench;